*** CIRCUITO RLC SÉRIE, GERADOR DE PULSO ALTA TENSÃO ***

C 1 0 0.6U IC=30E3V
R 1 2 11.56
L 2 0 108U

.end
