V1 5 0 2V
R1 5 1 100K
RF 3 1 500K
RP 2 0 1M
*AMPOP 
RI 2 1 1E12
RO 4 3 1M
EOP 4 0 2 1 1E10
*ENTRADA
Vdd 5 0 2V
.END

