R1 1 3 10K
R2 2 4 10K
R3 4 0 10K
R4 3 5 10K
R5 5 0 10K

*AMPOP 
RI 4 3 1E12
RO 6 5 1M
EOP 6 0 4 3 1E10

*ENTRADAS
Va1 1 0 3V
Va2 2 0 4V
.END

