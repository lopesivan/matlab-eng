BJT_DIFFAMP1.CIR - BJT DIFFERENTIAL AMPLIFIER
*
* SIGNAL SOURCE
VS	1	2	AC	1	SIN(0	10MVPEAK	10KHZ)
VCM	2	0	SIN(0	0MVPEAK	5KHZ)
*
* POWER SUPPLIES
VCC	11	0	DC	+15V
VDD	12	0	DC	-15V
*
Q1	3 1	5	Q2N2222
Q2	4 2	5	Q2N2222
RC1	11	3	1000
RC2	11	4	1000
RE	5	12	7.2K
*
*
.model Q2N2222  NPN(Is=3.108f Xti=3 Eg=1.11 Vaf=131.5 Bf=217.5 Ne=1.541
+               Ise=190.7f Ikf=1.296 Xtb=1.5 Br=6.18 Nc=2 Isc=0 Ikr=0 Rc=1
+               Cjc=14.57p Vjc=.75 Mjc=.3333 Fc=.5 Cje=26.08p Vje=.75
+               Mje=.3333 Tr=51.35n Tf=451p Itf=.1 Vtf=10 Xtf=2 Rb=10)
*
*
* CHECK DISTORTION WITH FOURIER SERIES ANALYSIS
.FOUR 10KHZ V(3,4)
*
* ANALYSIS
.TRAN 	5US  200US
.AC 	DEC 	5 1K 100MEG
*
* VIEW RESULTS
.PRINT	TRAN 	V(3) V(4)
.PRINT	AC 	V(3)
.PROBE
.END